----------------------------------------------------------------------------------
-- Company: Technical University of Cluj Napoca
-- Engineer: Chereja Iulia
-- Project Name: NAPOSIP
-- Description: Counter 74163 with activity monitoring 
--              - inputs:  CK, CLRN, LOADN, PT, D, C, B, A -std_logic  
--              - outputs : Qd, Qc, Qb, Qa, RCO -std_logic
--              - consumption :  port to monitor dynamic and static consumption
-- Dependencies: none
-- 
-- Revision: 1.0 - Added comments - Botond Sandor Kirei
-- Revision 0.01 - File Created
----------------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.std_logic_unsigned.all;

library work;
use work.PELib.all;
use work.PEGates.all;

entity num74163 is
    Generic (delay : time := 1 ns;
				 logic_family : logic_family_t; -- the logic family of the component
				 gate : component_t; -- the type of the component
				 Cload : real := 5.0 -- capacitive load 
                );
        Port ( CLK, CLRN, LOADN, P, T, D ,C ,B ,A : in std_logic;
                 Qd, Qc, Qb, Qa, RCO: out std_logic;
                 Vcc : in real ; -- supply voltage
		         consumption : out consumption_type := (0.0,0.0)
		         );
end num74163;

architecture Behavioral of num74163 is
signal counter : std_logic_vector (3 downto 0);
signal ck,cl,ld,en,dd,cc,bb,aa,qdd,qcc,qbb,qaa,rrco: std_logic;
begin
ck <= CLK;
cl <= CLRN;
ld <= LOADN;
en <= P;
dd <= D;
cc <= C;
bb <= B;
aa <= A;
functionare: process(ck,cl)
             begin
             if cl = '0' then
                   counter <= "0000";
             elsif rising_edge(ck) then
             if (ld = '0') then
                   counter <= dd & cc & bb & aa;
             elsif ( en = '1') then 
                   counter <= counter + 1;
       end if;
   end if;
end process;

qdd <= counter(3) after delay;
qcc <= counter(2) after delay;
qbb <= counter(1) after delay;
qaa <= counter(0) after delay;
rrco <= '1' after delay when (en = '1' and counter = "1111") else '0' after delay;

RCO <= rrco;
Qd <= qdd;
Qc <= qcc;
Qb <= qbb;
Qa <= qaa;

cm_i : consumption_monitor generic map ( N=>8, M=>5, logic_family => logic_family, gate => none_comp, Cload => Cload)
		port map (sin(0) => ck, sin(1) => cl, sin(2) => ld, sin(3) => en, sin(4) => dd, sin(5) => cc, sin(6) => bb, sin(7) => aa, Vcc => Vcc, sout(0) => qdd, sout(1) => qcc, sout(2) => qbb, sout(3) => qaa, sout(4) => rrco, consumption => consumption);
end Behavioral;


architecture Structural of num74163 is
-- implementation follows schematic in https://assets.nexperia.com/documents/data-sheet/74HC_HCT163.pdf
	signal CPn , MR, PE : std_logic;
	signal DFF0Qn, DFF1Qn, DFF2Qn, DFF3Qn : std_logic;
	signal DFF0Q, DFF1Q, DFF2Q, DFF3Q : std_logic;
	signal D0, D1, D2, D3 : std_logic;
	signal DFF0, DFF1, DFF2, DFF3 : std_logic;
	signal D01, D11, D21, D31 : std_logic;
	signal D02, D12, D22, D32 : std_logic;
	signal C0, C1, C2, C3 : std_logic;
	signal L0, L1, L2, L3, L31, L32 : std_logic;
	signal CET, CEP, TC, CE, Load, Reset : std_logic;
	signal net1, net2 : std_logic;
	signal cons : consumption_type_array(1 to 46);
begin

	dff0_I : dff generic map (delay => 1 ns, logic_family => logic_family, gate => none_comp) port map (CP => CPn, D => DFF0, RDn => '1', SDn => '1', Qn => DFF0Q, Q => DFF0Qn, Vcc => Vcc, consumption => cons(1));
	dff1_I : dff generic map (delay => 2 ns, logic_family => logic_family, gate => none_comp) port map (CP => CPn, D => DFF1, RDn => '1', SDn => '1', Qn => DFF1Q, Q => DFF1Qn, Vcc => Vcc, consumption => cons(2));
	dff2_I : dff generic map (delay => 1 ns, logic_family => logic_family, gate => none_comp) port map (CP => CPn, D => DFF2, RDn => '1', SDn => '1', Qn => DFF2Q, Q => DFF2Qn, Vcc => Vcc, consumption => cons(3));
	dff3_I : dff generic map (delay => 2 ns, logic_family => logic_family, gate => none_comp) port map (CP => CPn, D => DFF3, RDn => '1', SDn => '1', Qn => DFF3Q, Q => DFF3Qn, Vcc => Vcc,  consumption => cons(4));
	
	
	inv1: inv_gate generic map (delay => 0 ns, logic_family => logic_family, gate => inv_comp) port map (a => clk, Vcc => Vcc, y => CPn, consumption => cons(5));  --CPn <= not clk;
	inv2: inv_gate generic map (delay => 0 ns, logic_family => logic_family, gate => inv_comp) port map (a => DFF0Qn, Vcc => Vcc, y => Qa, consumption => cons(6));  --Qa <= not DFF0Qn;
	inv3: inv_gate generic map (delay => 0 ns, logic_family => logic_family, gate => inv_comp) port map (a => DFF1Qn, Vcc => Vcc, y => Qb, consumption => cons(7));  --Qb <= not DFF1Qn;
	inv4: inv_gate generic map (delay => 0 ns, logic_family => logic_family, gate => inv_comp) port map (a => DFF2Qn, Vcc => Vcc, y => Qc, consumption => cons(8)); --Qc <= not DFF2Qn;
	inv5: inv_gate generic map (delay => 0 ns, logic_family => logic_family, gate => inv_comp) port map (a => DFF3Qn, Vcc => Vcc, y => Qd, consumption => cons(9));--Qd <= not DFF3Qn;
	inv6: inv_gate generic map (delay => 0 ns, logic_family => logic_family, gate => inv_comp) port map (a => CLRN, Vcc => Vcc, y => MR, consumption => cons(10)); --MR <= not CLRN;
	
	tristate1: tristate_buf generic map (delay => 0 ns, logic_family => logic_family, gate => tristate_comp) port map (a => LOADN, en => '1',  Vcc => Vcc, y => PE, consumption => cons(11)); --PE <= LOADN;
	tristate2: tristate_buf generic map (delay => 0 ns, logic_family => logic_family, gate => tristate_comp) port map (a => A, en => '1',  Vcc => Vcc, y => D0, consumption => cons(12)); --D0 <= A; (--not A)
	tristate3: tristate_buf generic map (delay => 0 ns, logic_family => logic_family, gate => tristate_comp) port map (a => B, en => '1',  Vcc => Vcc, y => D1, consumption => cons(13));  --D1 <= B; (--not B)
	tristate4: tristate_buf generic map (delay => 0 ns, logic_family => logic_family, gate => tristate_comp) port map (a => C, en => '1',  Vcc => Vcc, y => D2, consumption => cons(14));  --D2 <= C; --not C;
	tristate5: tristate_buf generic map (delay => 0 ns, logic_family => logic_family, gate => tristate_comp) port map (a => D, en => '1',  Vcc => Vcc, y => D3, consumption => cons(15));  --D3 <= D; --not D;
	tristate6: tristate_buf generic map (delay => 0 ns, logic_family => logic_family, gate => tristate_comp) port map (a => T, en => '1',  Vcc => Vcc, y => CET, consumption => cons(16));  --CET <= T;
	tristate7: tristate_buf generic map (delay => 0 ns, logic_family => logic_family, gate => tristate_comp) port map (a => P, en => '1',  Vcc => Vcc, y => CEP, consumption => cons(17));  --CEP <= P;
	inv7: inv_gate generic map (delay => 0 ns, logic_family => logic_family, gate => inv_comp) port map (a => TC, Vcc => Vcc, y => RCO, consumption => cons(18));--RCO <= not TC;
	and5_gate1: and5_gate generic map (delay => 0 ns, logic_family => logic_family, gate => none_comp) port map ( a => DFF0Q, b => DFF1Q, c => DFF2Q, d => DFF3Q, e => CET, y => TC, Vcc => Vcc , consumption => cons(19)); --TC <= (DFF0Q and DFF1Q and DFF2Q and DFF3Q and CET);
	nand_gate1 : nand_gate generic map (delay => 0 ns, logic_family => logic_family, gate => nand_comp) port map (a => CET, b=> CEP, Vcc => Vcc, y => CE, consumption => cons(20)); --CE <=  CET nand CEP;
	
	nor_gate1: nor_gate generic map (delay => 0 ns, logic_family => logic_family, gate => nor_comp) port map (a => MR, b=> PE, Vcc => Vcc, y => LOAD, consumption => cons(21)); -- LOAD <= MR nor PE;
	nor_gate2: nor_gate generic map (delay => 0 ns, logic_family => logic_family, gate => nor_comp) port map (a => Load, b=> MR, Vcc => Vcc, y => Reset, consumption => cons(22)); --Reset <= Load nor MR;
	
	inv8: inv_gate generic map (delay => 0 ns, logic_family => logic_family, gate => inv_comp) port map (a => CE, Vcc => Vcc, y => C0, consumption => cons(23)); --C0 <= not CE;
	nor_gate3: nor_gate generic map (delay => 0 ns, logic_family => logic_family, gate => nor_comp) port map (a => CE, b=> DFF0Qn, Vcc => Vcc, y => C1, consumption => cons(24)); -- C1 <= CE nor DFF0Qn;
	or3_gate1: or3_gate generic map (delay => 0 ns, logic_family => logic_family, gate => none_comp) port map (a => CE, b=> DFF0Qn, c => DFF1Qn, Vcc => Vcc, y => net1, consumption => cons(25)); --(CE or DFF0Qn or DFF1Qn)
	inv9: inv_gate generic map (delay => 0 ns, logic_family => logic_family, gate => inv_comp) port map (a => net1, Vcc => Vcc, y => C2, consumption => cons(26));--	C2 <= not (CE or DFF0Qn or DFF1Qn);
    or4_gate1: or4_gate generic map (delay => 0 ns, logic_family => logic_family, gate => none_comp) port map (a => CE, b=> DFF0Qn, c => DFF1Qn, d => DFF2Qn, Vcc => Vcc, y => net2, consumption => cons(27)); --(CE or DFF0Qn or DFF1Qn or DFF2Qn)
    inv10: inv_gate generic map (delay => 0 ns, logic_family => logic_family, gate => inv_comp) port map (a => net2, Vcc => Vcc, y => C3, consumption => cons(28));--    C3 <= not (CE or DFF0Qn or DFF1Qn or DFF2Qn);
	
	xnor_gate1 : xnor_gate generic map (delay => 0 ns, logic_family => logic_family, gate => none_comp) port map (a => C0, b=> DFF0Qn, Vcc => Vcc, y => L0, consumption => cons(29)); --L0 <= C0 xnor DFF0Qn;
	xnor_gate2 : xnor_gate generic map (delay => 0 ns, logic_family => logic_family, gate => none_comp) port map (a => C1, b=> DFF1Qn, Vcc => Vcc, y => L1, consumption => cons(30));--L1 <= C1 xnor DFF1Qn;
	xnor_gate3 : xnor_gate generic map (delay => 0 ns, logic_family => logic_family, gate => none_comp) port map (a => C2, b=> DFF2Qn, Vcc => Vcc, y => L2, consumption => cons(31)); --L2 <= C2 xnor DFF2Qn;
	
	or_gate1: or_gate generic map (delay => 0 ns, logic_family => logic_family, gate => or_comp) port map (a => L31, b=> L32, Vcc => Vcc, y => L3, consumption => cons(32)); --L3 <= L31 or L32 (L3 <= C3 xnor DFF3Qn;)
    and_gate1: and_gate generic map (delay => 0 ns, logic_family => logic_family, gate => and_comp) port map (a => C3, b => DFF3Qn, Vcc => Vcc, y => L31, consumption => cons(33)); --L31 <= C3 and DFF3Qn;
    nor_gate4: nor_gate generic map (delay => 0 ns, logic_family => logic_family, gate => nor_comp) port map (a => C3, b => DFF3Qn, Vcc => Vcc, y => L32, consumption => cons(34)); --L32 <= C3 nor DFF3Qn;
    and_gate2: and_gate generic map (delay => 0 ns, logic_family => logic_family, gate => and_comp) port map (a => D0, b => load, Vcc => Vcc, y => D01, consumption => cons(35)); --D01 <= D0 and load;
    and_gate3: and_gate generic map (delay => 0 ns, logic_family => logic_family, gate => and_comp) port map (a => D1, b => load, Vcc => Vcc, y => D11, consumption => cons(36));--D11 <= D1 and load;
	and_gate4: and_gate generic map (delay => 0 ns, logic_family => logic_family, gate => and_comp) port map (a => D2, b => load, Vcc => Vcc, y => D21, consumption => cons(37));--D21 <= D2 and load;
	and_gate5: and_gate generic map (delay => 0 ns, logic_family => logic_family, gate => and_comp) port map (a => D3, b => load, Vcc => Vcc, y => D31, consumption => cons(38));--D31 <= D3 and load;
	and_gate6: and_gate generic map (delay => 0 ns, logic_family => logic_family, gate => and_comp) port map (a => L0, b => Reset, Vcc => Vcc, y => D02, consumption => cons(39)); --D02 <= L0 and Reset;
	and_gate7: and_gate generic map (delay => 0 ns, logic_family => logic_family, gate => and_comp) port map (a => L1, b=> Reset, Vcc => Vcc, y => D12, consumption => cons(40));--D12 <= L1 and Reset;
	and_gate8: and_gate generic map (delay => 0 ns, logic_family => logic_family, gate => and_comp) port map (a => L2, b=> Reset, Vcc => Vcc, y => D22, consumption => cons(41));--D22 <= L2 and Reset;
	and_gate9: and_gate generic map (delay => 0 ns, logic_family => logic_family, gate => and_comp) port map (a => L3, b=> Reset, Vcc => Vcc, y => D32, consumption => cons(42));--D32 <= L3 and Reset;
	
	nor_gate5: nor_gate generic map (delay => 0 ns, logic_family => logic_family, gate => nor_comp) port map (a => D01, b => D02, Vcc => Vcc, y => DFF0, consumption => cons(43));--DFF0 <= D01 nor D02;
	nor_gate6: nor_gate generic map (delay => 0 ns, logic_family => logic_family, gate => nor_comp) port map (a => D11, b => D12, Vcc => Vcc, y => DFF1, consumption => cons(44));--DFF1 <= D11 nor D12;
	nor_gate7: nor_gate generic map (delay => 0 ns, logic_family => logic_family, gate => nor_comp) port map (a => D21, b => D22, Vcc => Vcc, y => DFF2, consumption => cons(45));--DFF2 <= D21 nor D22;
	nor_gate8: nor_gate generic map (delay => 0 ns, logic_family => logic_family, gate => nor_comp) port map (a => D31, b => D32, Vcc => Vcc, y => DFF3, consumption => cons(46));--DFF3 <= D31 nor D32;
	
	sum : sum_up generic map (N => 46) port map (cons => cons, consumption => consumption );

	-- cm_i : consumption_monitor generic map (N=> 51, M => 5, Cin => Cin, Cpd => Cpd, Cload => Cload, Icc => Icc) port map (
	-- sin(0) => CPn	,
	-- sin(1) => DFF0Qn ,
	-- sin(2) => DFF1Qn ,
	-- sin(3) => DFF2Qn ,
	-- sin(4) => DFF3Qn ,
	-- sin(5) => DFF0Q  ,
	-- sin(6) => DFF1Q  ,
	-- sin(7) => DFF2Q  ,
	-- sin(8) => DFF3Q  ,
	-- sin(9) => MR     ,
	-- sin(10) => PE     ,
	-- sin(11) => D0     ,
	-- sin(12) => D1     ,
	-- sin(13) => D2     ,
	-- sin(14) => D3     ,
	-- sin(15) => CET    ,
	-- sin(16) => CEP    ,
	-- sin(17) => TC     ,
	-- sin(18) => CE     ,
	-- sin(19) => LOAD   ,
	-- sin(20) => Reset  ,
	-- sin(21) => C0     ,
	-- sin(22) => C1     ,
	-- sin(23) => C2     ,
	-- sin(24) => C3     ,
	-- sin(25) => L0     ,
	-- sin(26) => L1     ,
	-- sin(27) => L2     ,
	-- sin(28) => L3     ,
	-- sin(29) => L31    ,
	-- sin(30) => L32    ,
	-- sin(31) => D01    ,
	-- sin(32) => D11    ,
	-- sin(33) => D21    ,
	-- sin(34) => D31    ,
	-- sin(35) => D02    ,
	-- sin(36) => D12    ,
	-- sin(37) => D22    ,
	-- sin(38) => D32    ,
	-- sin(39) => DFF0   ,
	-- sin(40) => DFF1   ,
	-- sin(41) => DFF2   ,
	-- sin(42) => DFF3   ,
	-- sin(43) => CLK   ,
	-- sin(44) => CLRN  ,
	-- sin(45) => P ,
	-- sin(46) => T ,
	-- sin(47) => A ,
	-- sin(48) => B ,
	-- sin(49) => C ,
	-- sin(50) => D ,
	-- sout(0) => DFF0Qn , -- instead of Qa    ,
	-- sout(1) => DFF1Qn , -- instead of Qb    ,
	-- sout(2) => DFF2Qn , -- instead of Qc    ,
	-- sout(3) => DFF3Qn , -- instead of Qd    ,
	-- sout(4) => TC     , -- instead of RCO   ,
	-- consumption => cons(5));
	
	
end architecture;
